//------------------------------------------------------------------------------
// (c) ChipVerify
//------------------------------------------------------------------------------

module behave;
	reg [1:0]  a, b;

	initial begin
		a = 2'b10;
		#20  b = 2'b11;
	end

 	initial begin
		#10 a = 2'b11;
		#40 b = 2'b10;
	end

	initial 
		#60 $finish;
endmodule
